/*******************************************************
*  AN7   AN6   AN5   AN4  | AN3   AN2   AN1   AN0
*   |     |     |     |   |  |     |     |     |
*   __    __    __    __  |  __    __    __    __
*  |__|  |__|  |__|  |__| | |__|  |__|  |__|  |__|
*  |__|. |__|. |__|. |__|.| |__|. |__|. |__|. |__|.
*      
*  | |   | |   | |   | |  |  | |   | |   | |   | |
* CA CB CC CD CE CF CG DP | CA CB CC CD CE CF CG DP
********************************************************/

/********************************************************
*              _____
*          ___|  A  |___
*         |   |-----|   |
*         | F |     | B |
*         |___|-----|___|
*          ___|  G  |___
*         |   |-----|   |
*         | E |     | C |
*         |___|_____|___|     ---
*             |  D  |        | P |
*              -----          ---
*********************************************************/
module anode_control (
    input [2:0] refreshcounter,
    output reg [7:0] anode = 0
);

  always @(refreshcounter) begin
    case (refreshcounter)
      /*              |7|6|5|4|3|2|1|0|        */
      3'd0: anode = 8'b1_1_1_1_1_1_1_0;  // digit 1 ON
      3'd1: anode = 8'b1_1_1_1_1_1_0_1;  // digit 2 ON
      3'd2: anode = 8'b1_1_1_1_1_0_1_1;  // digit 3 ON
      3'd3: anode = 8'b1_1_1_1_0_1_1_1;  // digit 4 ON 
      3'd4: anode = 8'b1_1_1_0_1_1_1_1;  // digit 5 ON 
      3'd5: anode = 8'b1_1_1_1_1_1_1_1;  // digit 5 ON 
      3'd6: anode = 8'b1_1_1_1_1_1_1_1;  // digit 6 ON 
      3'd7: anode = 8'b0_1_1_1_1_1_1_1;  // digit 7 ON 
    endcase

  end

endmodule
